248503890f17ce512a2a07926841854a337bde567cfdf64500e64ab0
