077e7b8f9680b3260b7e5ccf22e8e7e701b79b195a5dfc4caa54cd6b
