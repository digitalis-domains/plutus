c89f700b5c7b8b060aba91e41ce31922f8742a6ac0b8865646ebfe90
